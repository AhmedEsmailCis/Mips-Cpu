----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    02:23:08 04/18/2018 
-- Design Name: 
-- Module Name:    mux2x1_32B - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity mux2x1_32B is
    Port ( R_type : in  STD_LOGIC_VECTOR (31 downto 0);
           I_type : in  STD_LOGIC_VECTOR (31 downto 0);
			   S : in  STD_LOGIC;
           ALU_data2 : out  STD_LOGIC_VECTOR (31 downto 0));
          
end mux2x1_32B;

architecture Behavioral of mux2x1_32B is

begin
ALU_data2<=R_type when S='0' else 
            I_type ;

end Behavioral;

